`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:54:11 01/15/2017 
// Design Name: 
// Module Name:    adder_8bits 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder_8bits(
	input  [7:0] in1,
	input  [7:0] in2,
	output [7:0] sum,
	output       c
	);


endmodule
